ENTITY detectacentena IS 
	PORT ( 	I1, I2, I3, I4, I5, I6 	: IN 	BIT ; 
		c : OUT 	BIT ) ; 
END detectacentena; 

ARCHITECTURE LogicFunc OF detectacentena IS 
BEGIN   

c <=
(I6 AND I5 AND (NOT I4) AND (NOT I3) AND I2 AND (NOT I1)) OR
(I6 AND I5 AND (NOT I4) AND (NOT I3) AND I2 AND I1) OR
(I6 AND I5 AND (NOT I4) AND I3 AND (NOT I2) AND (NOT I1)) OR
(I6 AND I5 AND (NOT I4) AND I3 AND (NOT I2) AND I1) OR
(I6 AND I5 AND (NOT I4) AND I3 AND I2 AND (NOT I1)) OR
(I6 AND I5 AND (NOT I4) AND I3 AND I2 AND I1) OR
(I6 AND I5 AND I4 AND (NOT I3) AND (NOT I2) AND (NOT I1)) OR
(I6 AND I5 AND I4 AND (NOT I3) AND (NOT I2) AND I1) OR
(I6 AND I5 AND I4 AND (NOT I3) AND I2 AND (NOT I1)) OR
(I6 AND I5 AND I4 AND (NOT I3) AND I2 AND I1) OR
(I6 AND I5 AND I4 AND I3 AND (NOT I2) AND (NOT I1)) OR
(I6 AND I5 AND I4 AND I3 AND (NOT I2) AND I1) OR
(I6 AND I5 AND I4 AND I3 AND I2 AND (NOT I1)) OR
(I6 AND I5 AND I4 AND I3 AND I2 AND I1);



END LogicFunc ;

