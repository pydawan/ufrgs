ENTITY conversorBin2Dec IS 
	PORT ( 	I1, I2, I3, I4, I5, I6 	: IN 	BIT ; 
		x2, x3, x4, y1, y2, y3, y4 : OUT 	BIT ) ; 
END conversorBin2Dec; 

ARCHITECTURE LogicFunc OF conversorBin2Dec IS 
BEGIN   
x2 <= 
((NOT I5 AND NOT I4 AND I3 AND I2 AND NOT I1)
OR
(NOT I6 AND NOT I5 AND I4 AND NOT I3 AND NOT I2 AND NOT I1)
OR
(NOT I6 AND NOT I5 AND I4 AND I3 AND NOT I2 AND I1)
OR
(NOT I6 AND I5 AND I4 AND I3 AND NOT I2 AND NOT I1)
OR
(I6 AND NOT I5 AND NOT I4 AND I3 AND NOT I1)
OR
(I6 AND NOT I5 AND I3 AND I2 AND NOT I1)
OR
(I6 AND I5 AND NOT I4 AND NOT I3 AND I2 AND I1)
OR
(NOT I6 AND NOT I5 AND NOT I4 AND NOT I3 AND I1)
OR
(I6 AND NOT I5 AND NOT I3 AND NOT I2 AND I1)
OR
(NOT I5 AND I4 AND NOT I3 AND I2 AND I1)
OR
(NOT I6 AND I5 AND NOT I4 AND NOT I3 AND NOT I1)
OR
(I6 AND I5 AND NOT I3 AND NOT I2 AND NOT I1)
OR
(I5 AND I4 AND NOT I3 AND I2 AND NOT I1)
OR
(I5 AND I4 AND I3 AND I2 AND I1)
OR
(NOT I6 AND I5 AND NOT I4 AND I3 AND I1)
OR
(I6 AND I5 AND I3 AND NOT I2 AND I1));

x3 <=
(((NOT I6) AND (NOT I5) AND I4 AND (NOT I2) AND (NOT I1)) OR
((NOT I6) AND (NOT I5) AND I4 AND I3 AND (NOT I2)) OR
((NOT I6) AND I5 AND (NOT I4) AND (NOT I3) AND (NOT I2) AND I1) OR
((NOT I6) AND I5 AND I4 AND (NOT I3) AND I2 AND I1) OR
((NOT I6) AND I4 AND I3 AND (NOT I2) AND (NOT I1)) OR
(I6 AND (NOT I5) AND (NOT I4) AND I3 AND I2 AND (NOT I1)) OR
(I6 AND I5 AND I4 AND (NOT I3) AND (NOT I2) AND I1) OR
((NOT I6) AND (NOT I5) AND (NOT I4) AND (NOT I3) AND I2) OR
((NOT I6) AND I5 AND (NOT I4) AND I2 AND (NOT I1)) OR
((NOT I6) AND (NOT I4) AND I3 AND I2 AND I1) OR
(I6 AND I5 AND I4 AND I2 AND (NOT I1)) OR
(I6 AND (NOT I5) AND I4 AND (NOT I3) AND I2) OR
(I6 AND I4 AND I3 AND I2 AND I1) OR
(I6 AND (NOT I5) AND (NOT I4) AND (NOT I3) AND (NOT I2)) OR
(I6 AND I5 AND (NOT I4) AND (NOT I2) AND (NOT I1)) OR
(I6 AND (NOT I4) AND I3 AND (NOT I2) AND I1));

x4 <=
(((NOT I6) AND (NOT I5)  AND (NOT I4) AND I3 AND (NOT I2)  AND (NOT I1) ) OR
((NOT I6) AND (NOT I5) AND I4 AND (NOT I3)  AND (NOT I2) AND I1) OR
((NOT I6) AND (NOT I5) AND I4 AND I3 AND I2 AND (NOT I1) ) OR
((NOT I6) AND I5 AND (NOT I4)  AND (NOT I3) AND I2 AND I1) OR
((NOT I6) AND I5 AND I4 AND (NOT I3)  AND (NOT I2)  AND (NOT I1) ) OR
((NOT I6) AND I5 AND I4 AND I3 AND (NOT I2) AND I1) OR
(I6 AND (NOT I5)  AND (NOT I4)  AND (NOT I3) AND I2 AND (NOT I1) ) OR
(I6 AND (NOT I5)  AND (NOT I4) AND I3 AND I2 AND I1) OR
(I6 AND (NOT I5) AND I4 AND I3 AND (NOT I2)  AND (NOT I1) ) OR
(I6 AND I5 AND (NOT I4)  AND (NOT I3)  AND (NOT I2) AND I1) OR
(I6 AND I5 AND (NOT I4) AND I3 AND I2 AND (NOT I1) ) OR
(I6 AND I5 AND I4 AND (NOT I3) AND I2 AND I1));

y1 <=
(((NOT I5)  AND (NOT I4) AND I3 AND I1) OR
((NOT I5)  AND (NOT I4) AND I3 AND I2) OR
((NOT I6) AND (NOT I5) AND I4 AND (NOT I3)  AND (NOT I2) ) OR
((NOT I5) AND I3 AND I2 AND I1) OR
((NOT I6) AND I5 AND I4 AND I3 AND (NOT I2) ) OR
(I6 AND (NOT I5)  AND (NOT I4) AND I2 AND I1) OR
(I6 AND (NOT I5)  AND (NOT I4) AND I3) OR
(I6 AND (NOT I5) AND I3 AND I1) OR
(I6 AND (NOT I5) AND I3 AND I2) OR
(I6 AND (NOT I4) AND I3 AND I2 AND I1) OR
(I5 AND (NOT I3)  AND (NOT I2) AND I1) OR
((NOT I6) AND I5 AND (NOT I3) AND I2) OR
(I6 AND I5 AND I4 AND (NOT I3) ) OR
(I5 AND (NOT I4)  AND (NOT I3)  AND (NOT I2)));

y2 <=
(((NOT I6) AND (NOT I5) AND I4 AND I2) OR
((NOT I6) AND (NOT I5) AND I4 AND I3) OR
((NOT I6) AND I5 AND (NOT I4) AND (NOT I3) ) OR
(I6 AND (NOT I5) AND (NOT I4) ) OR
(I6 AND I5 AND I4 AND I3) OR
((NOT I6) AND I4 AND I3 AND I2));

y3 <=
(((NOT I6) AND I5 AND I3) OR
((NOT I6) AND I5 AND I4) OR
(I6 AND (NOT I5) AND (NOT I4)));

y4 <=
((I6 AND (NOT I5) AND I4) OR
(I6 AND I5 AND (NOT I4) AND (NOT I3) AND (NOT I2)));



END LogicFunc ;

